module registerfile();
logic signed [63:0] gpr [31:0];
endmodule
