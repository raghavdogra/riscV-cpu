module registerfile();

logic signed [63:0] gpr [31:0];
logic signed  gprbusy [31:0];

endmodule
